`include"COM3to8Decoder";

module COM3to8Decoder_tb(
    reg [2:0] r;
    wire [7:0] w;
);

endmodule